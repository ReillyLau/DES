`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2018/04/11 19:59:08
// Design Name: 
// Module Name: key_sched
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module key_sched(
    input [63:0] key,
    output [47:0] subkey1,
    output [47:0] subkey2,
    output [47:0] subkey3,
    output [47:0] subkey4,
    output [47:0] subkey5,
    output [47:0] subkey6,
    output [47:0] subkey7,
    output [47:0] subkey8,
    output [47:0] subkey9,
    output [47:0] subkey10,
    output [47:0] subkey11,
    output [47:0] subkey12,
    output [47:0] subkey13,
    output [47:0] subkey14,
    output [47:0] subkey15,
    output [47:0] subkey16
    );

wire[55:0]		key_PC1;
wire[27:0]		c0, c1, c2, c3, c4, c5, c6, c7, c8, c9, c10, c11, c12, c13, c14, c15, c16;
wire[27:0]		d0, d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15, d16;

wire[55:0]		cd1, cd2, cd3, cd4, cd5, cd6, cd7, cd8, cd9, cd10, cd11, cd12, cd13, cd14, cd15, cd16;
/*************		初始密钥置换			*****************/
assign key_PC1 = {key[7], key[15], key[23], key[31], key[39], key[47], key[55], key[63], key[4], key[14], key[22], key[30], key[38], key[46], key[54], key[62], key[5], key[13], key[21], key[29], key[37], key[45], key[53], key[61], key[4], key[12], key[20], key[28], key[1], key[9], key[17], key[25], key[33], key[41], key[49], key[57], key[2], key[10], key[18], key[26], key[34], key[42], key[50], key[58], key[3], key[11], key[19], key[27], key[35], key[43], key[51], key[59], key[36], key[44], key[52], key[60]};

/****************	轮密钥置换			*************************/
assign subkey1 = {cd1[42], cd1[39], cd1[45], cd1[32], cd1[55], cd1[51], cd1[53], cd1[28], cd1[41], cd1[50], cd1[35], cd1[46], cd1[33], cd1[37], cd1[44], cd1[52], cd1[30], cd1[48], cd1[40], cd1[49], cd1[29], cd1[36], cd1[43], cd1[54], cd1[15], cd1[4], cd1[25], cd1[19], cd1[9], cd1[1], cd1[26], cd1[16], cd1[5], cd1[11], cd1[23], cd1[8], cd1[12], cd1[7], cd1[17], cd1[0], cd1[22], cd1[3], cd1[10], cd1[14], cd1[6], cd1[20], cd1[27], cd1[24]};

assign subkey2 = {cd2[42], cd2[39], cd2[45], cd2[32], cd2[55], cd2[51], cd2[53], cd2[28], cd2[41], cd2[50], cd2[35], cd2[46], cd2[33], cd2[37], cd2[44], cd2[52], cd2[30], cd2[48], cd2[40], cd2[49], cd2[29], cd2[36], cd2[43], cd2[54], cd2[15], cd2[4], cd2[25], cd2[19], cd2[9], cd2[1], cd2[26], cd2[16], cd2[5], cd2[11], cd2[23], cd2[8], cd2[12], cd2[7], cd2[17], cd2[0], cd2[22], cd2[3], cd2[10], cd2[14], cd2[6], cd2[20], cd2[27], cd2[24]};

assign subkey3 = {cd3[42], cd3[39], cd3[45], cd3[32], cd3[55], cd3[51], cd3[53], cd3[28], cd3[41], cd3[50], cd3[35], cd3[46], cd3[33], cd3[37], cd3[44], cd3[52], cd3[30], cd3[48], cd3[40], cd3[49], cd3[29], cd3[36], cd3[43], cd3[54], cd3[15], cd3[4], cd3[25], cd3[19], cd3[9], cd3[1], cd3[26], cd3[16], cd3[5], cd3[11], cd3[23], cd3[8], cd3[12], cd3[7], cd3[17], cd3[0], cd3[22], cd3[3], cd3[10], cd3[14], cd3[6], cd3[20], cd3[27], cd3[24]};

assign subkey4 = {cd4[42], cd4[39], cd4[45], cd4[32], cd4[55], cd4[51], cd4[53], cd4[28], cd4[41], cd4[50], cd4[35], cd4[46], cd4[33], cd4[37], cd4[44], cd4[52], cd4[30], cd4[48], cd4[40], cd4[49], cd4[29], cd4[36], cd4[43], cd4[54], cd4[15], cd4[4], cd4[25], cd4[19], cd4[9], cd4[1], cd4[26], cd4[16], cd4[5], cd4[11], cd4[23], cd4[8], cd4[12], cd4[7], cd4[17], cd4[0], cd4[22], cd4[3], cd4[10], cd4[14], cd4[6], cd4[20], cd4[27], cd4[24]};

assign subkey5 = {cd5[42], cd5[39], cd5[45], cd5[32], cd5[55], cd5[51], cd5[53], cd5[28], cd5[41], cd5[50], cd5[35], cd5[46], cd5[33], cd5[37], cd5[44], cd5[52], cd5[30], cd5[48], cd5[40], cd5[49], cd5[29], cd5[36], cd5[43], cd5[54], cd5[15], cd5[4], cd5[25], cd5[19], cd5[9], cd5[1], cd5[26], cd5[16], cd5[5], cd5[11], cd5[23], cd5[8], cd5[12], cd5[7], cd5[17], cd5[0], cd5[22], cd5[3], cd5[10], cd5[14], cd5[6], cd5[20], cd5[27], cd5[24]};

assign subkey6 = {cd6[42], cd6[39], cd6[45], cd6[32], cd6[55], cd6[51], cd6[53], cd6[28], cd6[41], cd6[50], cd6[35], cd6[46], cd6[33], cd6[37], cd6[44], cd6[52], cd6[30], cd6[48], cd6[40], cd6[49], cd6[29], cd6[36], cd6[43], cd6[54], cd6[15], cd6[4], cd6[25], cd6[19], cd6[9], cd6[1], cd6[26], cd6[16], cd6[5], cd6[11], cd6[23], cd6[8], cd6[12], cd6[7], cd6[17], cd6[0], cd6[22], cd6[3], cd6[10], cd6[14], cd6[6], cd6[20], cd6[27], cd6[24]};

assign subkey7 = {cd7[42], cd7[39], cd7[45], cd7[32], cd7[55], cd7[51], cd7[53], cd7[28], cd7[41], cd7[50], cd7[35], cd7[46], cd7[33], cd7[37], cd7[44], cd7[52], cd7[30], cd7[48], cd7[40], cd7[49], cd7[29], cd7[36], cd7[43], cd7[54], cd7[15], cd7[4], cd7[25], cd7[19], cd7[9], cd7[1], cd7[26], cd7[16], cd7[5], cd7[11], cd7[23], cd7[8], cd7[12], cd7[7], cd7[17], cd7[0], cd7[22], cd7[3], cd7[10], cd7[14], cd7[6], cd7[20], cd7[27], cd7[24]};

assign subkey8 = {cd8[42], cd8[39], cd8[45], cd8[32], cd8[55], cd8[51], cd8[53], cd8[28], cd8[41], cd8[50], cd8[35], cd8[46], cd8[33], cd8[37], cd8[44], cd8[52], cd8[30], cd8[48], cd8[40], cd8[49], cd8[29], cd8[36], cd8[43], cd8[54], cd8[15], cd8[4], cd8[25], cd8[19], cd8[9], cd8[1], cd8[26], cd8[16], cd8[5], cd8[11], cd8[23], cd8[8], cd8[12], cd8[7], cd8[17], cd8[0], cd8[22], cd8[3], cd8[10], cd8[14], cd8[6], cd8[20], cd8[27], cd8[24]};

assign subkey9 = {cd9[42], cd9[39], cd9[45], cd9[32], cd9[55], cd9[51], cd9[53], cd9[28], cd9[41], cd9[50], cd9[35], cd9[46], cd9[33], cd9[37], cd9[44], cd9[52], cd9[30], cd9[48], cd9[40], cd9[49], cd9[29], cd9[36], cd9[43], cd9[54], cd9[15], cd9[4], cd9[25], cd9[19], cd9[9], cd9[1], cd9[26], cd9[16], cd9[5], cd9[11], cd9[23], cd9[8], cd9[12], cd9[7], cd9[17], cd9[0], cd9[22], cd9[3], cd9[10], cd9[14], cd9[6], cd9[20], cd9[27], cd9[24]};

assign subkey10 = {cd10[42], cd10[39], cd10[45], cd10[32], cd10[55], cd10[51], cd10[53], cd10[28], cd10[41], cd10[50], cd10[35], cd10[46], cd10[33], cd10[37], cd10[44], cd10[52], cd10[30], cd10[48], cd10[40], cd10[49], cd10[29], cd10[36], cd10[43], cd10[54], cd10[15], cd10[4], cd10[25], cd10[19], cd10[9], cd10[1], cd10[26], cd10[16], cd10[5], cd10[11], cd10[23], cd10[8], cd10[12], cd10[7], cd10[17], cd10[0], cd10[22], cd10[3], cd10[10], cd10[14], cd10[6], cd10[20], cd10[27], cd10[24]};

assign subkey11 = {cd11[42], cd11[39], cd11[45], cd11[32], cd11[55], cd11[51], cd11[53], cd11[28], cd11[41], cd11[50], cd11[35], cd11[46], cd11[33], cd11[37], cd11[44], cd11[52], cd11[30], cd11[48], cd11[40], cd11[49], cd11[29], cd11[36], cd11[43], cd11[54], cd11[15], cd11[4], cd11[25], cd11[19], cd11[9], cd11[1], cd11[26], cd11[16], cd11[5], cd11[11], cd11[23], cd11[8], cd11[12], cd11[7], cd11[17], cd11[0], cd11[22], cd11[3], cd11[10], cd11[14], cd11[6], cd11[20], cd11[27], cd11[24]};

assign subkey12 = {cd12[42], cd12[39], cd12[45], cd12[32], cd12[55], cd12[51], cd12[53], cd12[28], cd12[41], cd12[50], cd12[35], cd12[46], cd12[33], cd12[37], cd12[44], cd12[52], cd12[30], cd12[48], cd12[40], cd12[49], cd12[29], cd12[36], cd12[43], cd12[54], cd12[15], cd12[4], cd12[25], cd12[19], cd12[9], cd12[1], cd12[26], cd12[16], cd12[5], cd12[11], cd12[23], cd12[8], cd12[12], cd12[7], cd12[17], cd12[0], cd12[22], cd12[3], cd12[10], cd12[14], cd12[6], cd12[20], cd12[27], cd12[24]};

assign subkey13 = {cd13[42], cd13[39], cd13[45], cd13[32], cd13[55], cd13[51], cd13[53], cd13[28], cd13[41], cd13[50], cd13[35], cd13[46], cd13[33], cd13[37], cd13[44], cd13[52], cd13[30], cd13[48], cd13[40], cd13[49], cd13[29], cd13[36], cd13[43], cd13[54], cd13[15], cd13[4], cd13[25], cd13[19], cd13[9], cd13[1], cd13[26], cd13[16], cd13[5], cd13[11], cd13[23], cd13[8], cd13[12], cd13[7], cd13[17], cd13[0], cd13[22], cd13[3], cd13[10], cd13[14], cd13[6], cd13[20], cd13[27], cd13[24]};

assign subkey14 = {cd14[42], cd14[39], cd14[45], cd14[32], cd14[55], cd14[51], cd14[53], cd14[28], cd14[41], cd14[50], cd14[35], cd14[46], cd14[33], cd14[37], cd14[44], cd14[52], cd14[30], cd14[48], cd14[40], cd14[49], cd14[29], cd14[36], cd14[43], cd14[54], cd14[15], cd14[4], cd14[25], cd14[19], cd14[9], cd14[1], cd14[26], cd14[16], cd14[5], cd14[11], cd14[23], cd14[8], cd14[12], cd14[7], cd14[17], cd14[0], cd14[22], cd14[3], cd14[10], cd14[14], cd14[6], cd14[20], cd14[27], cd14[24]};

assign subkey15 = {cd15[42], cd15[39], cd15[45], cd15[32], cd15[55], cd15[51], cd15[53], cd15[28], cd15[41], cd15[50], cd15[35], cd15[46], cd15[33], cd15[37], cd15[44], cd15[52], cd15[30], cd15[48], cd15[40], cd15[49], cd15[29], cd15[36], cd15[43], cd15[54], cd15[15], cd15[4], cd15[25], cd15[19], cd15[9], cd15[1], cd15[26], cd15[16], cd15[5], cd15[11], cd15[23], cd15[8], cd15[12], cd15[7], cd15[17], cd15[0], cd15[22], cd15[3], cd15[10], cd15[14], cd15[6], cd15[20], cd15[27], cd15[24]};

assign subkey16 = {cd16[42], cd16[39], cd16[45], cd16[32], cd16[55], cd16[51], cd16[53], cd16[28], cd16[41], cd16[50], cd16[35], cd16[46], cd16[33], cd16[37], cd16[44], cd16[52], cd16[30], cd16[48], cd16[40], cd16[49], cd16[29], cd16[36], cd16[43], cd16[54], cd16[15], cd16[4], cd16[25], cd16[19], cd16[9], cd16[1], cd16[26], cd16[16], cd16[5], cd16[11], cd16[23], cd16[8], cd16[12], cd16[7], cd16[17], cd16[0], cd16[22], cd16[3], cd16[10], cd16[14], cd16[6], cd16[20], cd16[27], cd16[24]};

/*********		产生子密钥				*******************/
assign c0 = key_PC1[55:28];
assign d0 = key_PC1[27:0];
//
assign c1 = {c0[26:0], c0[27]};
assign d1 = {d0[26:0], d0[27]};
assign cd1 = {c1, d1};
//
assign c2 = {c1[26:0], c1[27]};
assign d2 = {d1[26:0], d1[27]};
assign cd2 = {c2, d2};
//
assign c3 = {c2[25:0], c2[27:26]};
assign d3 = {d2[25:0], d2[27:26]};
assign cd3 = {c3, d3};
//
assign c4 = {c3[25:0], c3[27:26]};
assign d4 = {d3[25:0], d3[27:26]};
assign cd4 = {c4, d4};
//
assign c5 = {c4[25:0], c4[27:26]};
assign d5 = {d4[25:0], d4[27:26]};
assign cd5 = {c5, d5};
//
assign c6 = {c5[25:0], c5[27:26]};
assign d6 = {d5[25:0], d5[27:26]};
assign cd6 = {c6, d6};
//
assign c7 = {c6[25:0], c6[27:26]};
assign d7 = {d6[25:0], d6[27:26]};
assign cd7 = {c7, d7};
//
assign c8 = {c7[25:0], c7[27:26]};
assign d8 = {d7[25:0], d7[27:26]};
assign cd8 = {c8, d8};
//
assign c9 = {c8[26:0], c8[27]};
assign d9 = {d8[26:0], d8[27]};
assign cd9 = {c9, d9};
//
assign c10 = {c9[25:0], c9[27:26]};
assign d10 = {d9[25:0], d9[27:26]};
assign cd10 = {c10, d10};
//
assign c11 = {c10[25:0], c10[27:26]};
assign d11 = {d10[25:0], d10[27:26]};
assign cd11 = {c11, d11};
//
assign c12 = {c11[25:0], c11[27:26]};
assign d12 = {d11[25:0], d11[27:26]};
assign cd12 = {c12, d12};
//
assign c13 = {c12[25:0], c12[27:26]};
assign d13 = {d12[25:0], d12[27:26]};
assign cd13 = {c13, d13};
//
assign c14 = {c13[25:0], c13[27:26]};
assign d14 = {d13[25:0], d13[27:26]};
assign cd14 = {c14, d14};
//
assign c15 = {c14[25:0], c14[27:26]};
assign d15 = {d14[25:0], d14[27:26]};
assign cd15 = {c15, d15};
//
assign c16 = {c15[26:0], c15[27]};
assign d16 = {d15[26:0], d15[27]};
assign cd16 = {c16, d16};
	
	
	
endmodule
